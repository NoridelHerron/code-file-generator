
// ===========================================================
// Project Name: 
// Description :
//
// File Name   : vc.v
// Dependencies:
// Author      : kjskjdsa
// Date        : 2026-01-09 10:46:37
// ===========================================================

module vc (
    
        // User/s
        // I/O
        
);

// Add wire or reg here


always @(*) begin
    // logic here
end

