
// ============================================================
// Project Name: 
// Description :
//
// File Name   : verilog_test.v
// Dependencies:
// Author      : Noriddel
// Date        : 2026-01-10 09:12:21
// ============================================================
`timescale 1ns / 1ps

module verilog_test (
    
        // User/s
        // I/O
        
);

// Add wire or reg here

always @(*) begin
    // logic here
end

