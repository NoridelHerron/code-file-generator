
// ============================================================
// Project Name: 
// Description :
//
// File Name   : verilog.vh
// Dependencies:
// Author      : sdfkjjs
// Date        : 2026-01-10 09:26:00
// ============================================================

`ifndef VERILOG_VH
`define VERILOG_VH

// parameters
// `define MACROS
// localparams

`endif

