
// ============================================================
// Project Name: 
// Description :
//
// File Name   : svh.svh
// Dependencies:
// Author      : Noridel
// Date        : 2026-01-10 17:05:51
// ============================================================

package svh_pkg;

    // parameters
    // typedefs
    // localparams
    // functions

endpackage

============================================================
// End of File
============================================================

