
-- ============================================================
-- Project Name: 
-- Description :
--
-- File Name   : vhdl.vhd
-- Dependencies:
-- Author      : jksa
-- Date        : 2026-01-10 17:54:45
-- ============================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- CUSTOMIZED PACKAGE
-- library work;
-- use work.xxxxxxx.all;

package vhdl_pkg is

    -- constants
    -- types
    -- subtypes
    -- function/procedure declarations

end package vhdl_pkg;

-- ****************************************

package body vhdl_pkg is

    -- function/procedure implementations

end package body vhdl_pkg;

-- ============================================================
-- END OF FILE
-- ============================================================

