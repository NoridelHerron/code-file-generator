
// ============================================================
// Project Name: 
// Description :
//
// File Name   : sv.svh
// Dependencies:
// Author      : kljdsfks
// Date        : 2026-01-10 09:26:45
// ============================================================

package sv_pkg;

    // parameters
    // typedefs
    // localparams
    // functions

endpackage

============================================================
// End of File
============================================================

