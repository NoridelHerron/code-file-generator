
// ===========================================================
// Project Name: 
// Description :
//
// File Name   : svc.sv
// Dependencies:
// Author      : Noride
// Date        : 2026-01-09 11:12:01
// ===========================================================

module svc (
    
        // User/s
        // I/O
        
);

// Add logic signal/s here


always_comb begin
    // logic here
end
    
