
// ===========================================================
// Project Name: 
// Description :
//
// File Name   : vh_pkg.vh
// Dependencies:
// Author      : Nor
// Date        : 2026-01-09 11:07:57
// ===========================================================

`ifndef VH_VH
`define VH_VH

// parameters
// `define MACROS
// localparams

`endif

