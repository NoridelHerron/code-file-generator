-- ============================================================
-- Project Name: 
-- Description :
--
-- File Name   : vhdl_c.vhd
-- Dependencies:
-- Author      : ajdh
-- Date        : 2026-01-10 19:15:59
-- ============================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- CUSTOMIZED PACKAGE
-- library work;
-- use work.xxxxxxx.all;

entity vhdl_c is
    port (

        -- User/s
        -- add ports here
        
    );
end vhdl_c;

architecture rtl of vhdl_c is

begin

    -- Combinational logic
    -- If only simple concurrent assignments are needed,
    -- this process can be safely removed.
    process(all)
    begin
        -- logic here
    end process;
    
end rtl;

-- ============================================================
-- END OF FILE
-- ============================================================
