
// ===========================================================
// Project Name: 
// Description :
//
// File Name   : v_test_pkg.vh
// Dependencies:
// Author      : Njkafjdf hdafhjhafh
// Date        : 2026-01-07 22:23:08
// ===========================================================

`ifndef V_TEST_PKG_VH
`define V_TEST_PKG_VH

// parameters
// `define MACROS
// localparams

`endif

