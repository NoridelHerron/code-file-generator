
// ============================================================
// Project Name: 
// Description :
//
// File Name   : vh.vh
// Dependencies:
// Author      : Nor
// Date        : 2026-01-10 17:06:29
// ============================================================

`ifndef VH_VH
`define VH_VH

// parameters
// `define MACROS
// localparams

`endif

