
// ============================================================
// Project Name: 
// Description :
//
// File Name   : svh.svh
// Dependencies:
// Author      : kjasd
// Date        : 2026-01-10 18:06:10
// ============================================================

package svh_pkg;

    // parameters
    // typedefs
    // localparams
    // functions

endpackage

// ============================================================
// End of File
// ============================================================

