
// ===========================================================
// Project Name: 
// Description :
//
// File Name   : sv_test_pkg.svh
// Dependencies:
// Author      : Nsooo
// Date        : 2026-01-07 22:24:52
// ===========================================================

package sv_test_pkg;

    // parameters
    // typedefs
    // localparams
    // functions

endpackage

