
// ===========================================================
// Project Name: 
// Description :
//
// File Name   : svh_pkg.svh
// Dependencies:
// Author      : jkldaj avjkjkd akjfjdf
// Date        : 2026-01-09 11:13:33
// ===========================================================

package svh;

    // parameters
    // typedefs
    // localparams
    // functions

endpackage

